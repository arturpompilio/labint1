// SistemaEmbarcado.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SistemaEmbarcado (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         conduit_img_1_done_write;                                    // Conduit_Img_1:done -> Subtrator:done1
	wire         conduit_img_2_done_write;                                    // Conduit_Img_2:done -> Subtrator:done2
	wire  [31:0] conduit_img_1_pixel_readdata;                                // Conduit_Img_1:read_conduit -> Subtrator:writedata1
	wire  [31:0] conduit_img_2_pixel_readdata;                                // Conduit_Img_2:read_conduit -> Subtrator:writedata2
	wire  [31:0] processador_data_master_readdata;                            // mm_interconnect_0:Processador_data_master_readdata -> Processador:d_readdata
	wire         processador_data_master_waitrequest;                         // mm_interconnect_0:Processador_data_master_waitrequest -> Processador:d_waitrequest
	wire         processador_data_master_debugaccess;                         // Processador:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Processador_data_master_debugaccess
	wire  [18:0] processador_data_master_address;                             // Processador:d_address -> mm_interconnect_0:Processador_data_master_address
	wire   [3:0] processador_data_master_byteenable;                          // Processador:d_byteenable -> mm_interconnect_0:Processador_data_master_byteenable
	wire         processador_data_master_read;                                // Processador:d_read -> mm_interconnect_0:Processador_data_master_read
	wire         processador_data_master_write;                               // Processador:d_write -> mm_interconnect_0:Processador_data_master_write
	wire  [31:0] processador_data_master_writedata;                           // Processador:d_writedata -> mm_interconnect_0:Processador_data_master_writedata
	wire  [31:0] processador_instruction_master_readdata;                     // mm_interconnect_0:Processador_instruction_master_readdata -> Processador:i_readdata
	wire         processador_instruction_master_waitrequest;                  // mm_interconnect_0:Processador_instruction_master_waitrequest -> Processador:i_waitrequest
	wire  [16:0] processador_instruction_master_address;                      // Processador:i_address -> mm_interconnect_0:Processador_instruction_master_address
	wire         processador_instruction_master_read;                         // Processador:i_read -> mm_interconnect_0:Processador_instruction_master_read
	wire         mm_interconnect_0_medidor_escrita_write;                     // mm_interconnect_0:Medidor_Escrita_write -> Medidor:write
	wire  [31:0] mm_interconnect_0_medidor_escrita_writedata;                 // mm_interconnect_0:Medidor_Escrita_writedata -> Medidor:writedata
	wire         mm_interconnect_0_conduit_img_1_escrita_write;               // mm_interconnect_0:Conduit_Img_1_Escrita_write -> Conduit_Img_1:write
	wire  [31:0] mm_interconnect_0_conduit_img_1_escrita_writedata;           // mm_interconnect_0:Conduit_Img_1_Escrita_writedata -> Conduit_Img_1:writedata
	wire         mm_interconnect_0_conduit_img_2_escrita_write;               // mm_interconnect_0:Conduit_Img_2_Escrita_write -> Conduit_Img_2:write
	wire  [31:0] mm_interconnect_0_conduit_img_2_escrita_writedata;           // mm_interconnect_0:Conduit_Img_2_Escrita_writedata -> Conduit_Img_2:writedata
	wire  [31:0] mm_interconnect_0_medidor_leitura_readdata;                  // Medidor:readdata -> mm_interconnect_0:Medidor_Leitura_readdata
	wire         mm_interconnect_0_medidor_leitura_read;                      // mm_interconnect_0:Medidor_Leitura_read -> Medidor:read
	wire  [31:0] mm_interconnect_0_conduit_img_1_leitura_readdata;            // Conduit_Img_1:readdata -> mm_interconnect_0:Conduit_Img_1_Leitura_readdata
	wire         mm_interconnect_0_conduit_img_1_leitura_read;                // mm_interconnect_0:Conduit_Img_1_Leitura_read -> Conduit_Img_1:read
	wire  [31:0] mm_interconnect_0_conduit_img_2_leitura_readdata;            // Conduit_Img_2:readdata -> mm_interconnect_0:Conduit_Img_2_Leitura_readdata
	wire         mm_interconnect_0_conduit_img_2_leitura_read;                // mm_interconnect_0:Conduit_Img_2_Leitura_read -> Conduit_Img_2:read
	wire  [31:0] mm_interconnect_0_subtrator_leitura_readdata;                // Subtrator:readdata -> mm_interconnect_0:Subtrator_Leitura_readdata
	wire         mm_interconnect_0_subtrator_leitura_read;                    // mm_interconnect_0:Subtrator_Leitura_read -> Subtrator:read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_processador_debug_mem_slave_readdata;      // Processador:debug_mem_slave_readdata -> mm_interconnect_0:Processador_debug_mem_slave_readdata
	wire         mm_interconnect_0_processador_debug_mem_slave_waitrequest;   // Processador:debug_mem_slave_waitrequest -> mm_interconnect_0:Processador_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_processador_debug_mem_slave_debugaccess;   // mm_interconnect_0:Processador_debug_mem_slave_debugaccess -> Processador:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_processador_debug_mem_slave_address;       // mm_interconnect_0:Processador_debug_mem_slave_address -> Processador:debug_mem_slave_address
	wire         mm_interconnect_0_processador_debug_mem_slave_read;          // mm_interconnect_0:Processador_debug_mem_slave_read -> Processador:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_processador_debug_mem_slave_byteenable;    // mm_interconnect_0:Processador_debug_mem_slave_byteenable -> Processador:debug_mem_slave_byteenable
	wire         mm_interconnect_0_processador_debug_mem_slave_write;         // mm_interconnect_0:Processador_debug_mem_slave_write -> Processador:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_processador_debug_mem_slave_writedata;     // mm_interconnect_0:Processador_debug_mem_slave_writedata -> Processador:debug_mem_slave_writedata
	wire         mm_interconnect_0_memoriaprograma_s1_chipselect;             // mm_interconnect_0:MemoriaPrograma_s1_chipselect -> MemoriaPrograma:chipselect
	wire  [31:0] mm_interconnect_0_memoriaprograma_s1_readdata;               // MemoriaPrograma:readdata -> mm_interconnect_0:MemoriaPrograma_s1_readdata
	wire  [13:0] mm_interconnect_0_memoriaprograma_s1_address;                // mm_interconnect_0:MemoriaPrograma_s1_address -> MemoriaPrograma:address
	wire   [3:0] mm_interconnect_0_memoriaprograma_s1_byteenable;             // mm_interconnect_0:MemoriaPrograma_s1_byteenable -> MemoriaPrograma:byteenable
	wire         mm_interconnect_0_memoriaprograma_s1_write;                  // mm_interconnect_0:MemoriaPrograma_s1_write -> MemoriaPrograma:write
	wire  [31:0] mm_interconnect_0_memoriaprograma_s1_writedata;              // mm_interconnect_0:MemoriaPrograma_s1_writedata -> MemoriaPrograma:writedata
	wire         mm_interconnect_0_memoriaprograma_s1_clken;                  // mm_interconnect_0:MemoriaPrograma_s1_clken -> MemoriaPrograma:clken
	wire         mm_interconnect_0_memoriaimg1_s1_chipselect;                 // mm_interconnect_0:MemoriaImg1_s1_chipselect -> MemoriaImg1:chipselect
	wire   [7:0] mm_interconnect_0_memoriaimg1_s1_readdata;                   // MemoriaImg1:readdata -> mm_interconnect_0:MemoriaImg1_s1_readdata
	wire         mm_interconnect_0_memoriaimg1_s1_debugaccess;                // mm_interconnect_0:MemoriaImg1_s1_debugaccess -> MemoriaImg1:debugaccess
	wire  [16:0] mm_interconnect_0_memoriaimg1_s1_address;                    // mm_interconnect_0:MemoriaImg1_s1_address -> MemoriaImg1:address
	wire         mm_interconnect_0_memoriaimg1_s1_write;                      // mm_interconnect_0:MemoriaImg1_s1_write -> MemoriaImg1:write
	wire   [7:0] mm_interconnect_0_memoriaimg1_s1_writedata;                  // mm_interconnect_0:MemoriaImg1_s1_writedata -> MemoriaImg1:writedata
	wire         mm_interconnect_0_memoriaimg1_s1_clken;                      // mm_interconnect_0:MemoriaImg1_s1_clken -> MemoriaImg1:clken
	wire         mm_interconnect_0_memoriaimg2_s1_chipselect;                 // mm_interconnect_0:MemoriaImg2_s1_chipselect -> MemoriaImg2:chipselect
	wire   [7:0] mm_interconnect_0_memoriaimg2_s1_readdata;                   // MemoriaImg2:readdata -> mm_interconnect_0:MemoriaImg2_s1_readdata
	wire         mm_interconnect_0_memoriaimg2_s1_debugaccess;                // mm_interconnect_0:MemoriaImg2_s1_debugaccess -> MemoriaImg2:debugaccess
	wire  [16:0] mm_interconnect_0_memoriaimg2_s1_address;                    // mm_interconnect_0:MemoriaImg2_s1_address -> MemoriaImg2:address
	wire         mm_interconnect_0_memoriaimg2_s1_write;                      // mm_interconnect_0:MemoriaImg2_s1_write -> MemoriaImg2:write
	wire   [7:0] mm_interconnect_0_memoriaimg2_s1_writedata;                  // mm_interconnect_0:MemoriaImg2_s1_writedata -> MemoriaImg2:writedata
	wire         mm_interconnect_0_memoriaimg2_s1_clken;                      // mm_interconnect_0:MemoriaImg2_s1_clken -> MemoriaImg2:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] processador_irq_irq;                                         // irq_mapper:sender_irq -> Processador:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Conduit_Img_1:reset_n, Conduit_Img_2:reset_n, Medidor:reset_n, MemoriaImg1:reset, MemoriaImg2:reset, MemoriaPrograma:reset, Processador:reset_n, Subtrator:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:Processador_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [MemoriaImg1:reset_req, MemoriaImg2:reset_req, MemoriaPrograma:reset_req, Processador:reset_req, rst_translator:reset_req_in]
	wire         processador_debug_reset_request_reset;                       // Processador:debug_reset_request -> rst_controller:reset_in1

	Reader_Interface conduit_img_1 (
		.clk          (clk_clk),                                           //   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                   //   reset.reset_n
		.readdata     (mm_interconnect_0_conduit_img_1_leitura_readdata),  // Leitura.readdata
		.read         (mm_interconnect_0_conduit_img_1_leitura_read),      //        .read
		.write        (mm_interconnect_0_conduit_img_1_escrita_write),     // Escrita.write
		.writedata    (mm_interconnect_0_conduit_img_1_escrita_writedata), //        .writedata
		.done         (conduit_img_1_done_write),                          //    Done.write
		.read_conduit (conduit_img_1_pixel_readdata)                       //   Pixel.readdata
	);

	Reader_Interface conduit_img_2 (
		.clk          (clk_clk),                                           //   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                   //   reset.reset_n
		.readdata     (mm_interconnect_0_conduit_img_2_leitura_readdata),  // Leitura.readdata
		.read         (mm_interconnect_0_conduit_img_2_leitura_read),      //        .read
		.write        (mm_interconnect_0_conduit_img_2_escrita_write),     // Escrita.write
		.writedata    (mm_interconnect_0_conduit_img_2_escrita_writedata), //        .writedata
		.done         (conduit_img_2_done_write),                          //    Done.write
		.read_conduit (conduit_img_2_pixel_readdata)                       //   Pixel.readdata
	);

	Clock_Counter_Interface medidor (
		.clk       (clk_clk),                                     //   clock.clk
		.reset_n   (~rst_controller_reset_out_reset),             //   reset.reset_n
		.write     (mm_interconnect_0_medidor_escrita_write),     // Escrita.write
		.writedata (mm_interconnect_0_medidor_escrita_writedata), //        .writedata
		.read      (mm_interconnect_0_medidor_leitura_read),      // Leitura.read
		.readdata  (mm_interconnect_0_medidor_leitura_readdata)   //        .readdata
	);

	SistemaEmbarcado_MemoriaImg1 memoriaimg1 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_memoriaimg1_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_memoriaimg1_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_memoriaimg1_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_memoriaimg1_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_memoriaimg1_s1_write),       //       .write
		.readdata    (mm_interconnect_0_memoriaimg1_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_memoriaimg1_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	SistemaEmbarcado_MemoriaImg2 memoriaimg2 (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_memoriaimg2_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_memoriaimg2_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_memoriaimg2_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_memoriaimg2_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_memoriaimg2_s1_write),       //       .write
		.readdata    (mm_interconnect_0_memoriaimg2_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_memoriaimg2_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	SistemaEmbarcado_MemoriaPrograma memoriaprograma (
		.clk        (clk_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_memoriaprograma_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoriaprograma_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoriaprograma_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoriaprograma_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoriaprograma_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoriaprograma_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoriaprograma_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),              //       .reset_req
		.freeze     (1'b0)                                             // (terminated)
	);

	SistemaEmbarcado_Processador processador (
		.clk                                 (clk_clk),                                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                           //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                           (processador_data_master_address),                           //               data_master.address
		.d_byteenable                        (processador_data_master_byteenable),                        //                          .byteenable
		.d_read                              (processador_data_master_read),                              //                          .read
		.d_readdata                          (processador_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (processador_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (processador_data_master_write),                             //                          .write
		.d_writedata                         (processador_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (processador_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (processador_instruction_master_address),                    //        instruction_master.address
		.i_read                              (processador_instruction_master_read),                       //                          .read
		.i_readdata                          (processador_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (processador_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (processador_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (processador_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_processador_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_processador_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_processador_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_processador_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_processador_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_processador_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_processador_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_processador_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                           // custom_instruction_master.readra
	);

	Teste_Subtrator_Interface subtrator (
		.clk        (clk_clk),                                      //       clock.clk
		.reset_n    (~rst_controller_reset_out_reset),              //       reset.reset_n
		.read       (mm_interconnect_0_subtrator_leitura_read),     //     Leitura.read
		.readdata   (mm_interconnect_0_subtrator_leitura_readdata), //            .readdata
		.writedata1 (conduit_img_1_pixel_readdata),                 // Pixel_Img_1.readdata
		.writedata2 (conduit_img_2_pixel_readdata),                 // Pixel_Img_2.readdata
		.done1      (conduit_img_1_done_write),                     //   Done_Img1.write
		.done2      (conduit_img_2_done_write)                      //   Done_Img2.write
	);

	SistemaEmbarcado_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	SistemaEmbarcado_mm_interconnect_0 mm_interconnect_0 (
		.Clock_clk_clk                                 (clk_clk),                                                     //                               Clock_clk.clk
		.Processador_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // Processador_reset_reset_bridge_in_reset.reset
		.Processador_data_master_address               (processador_data_master_address),                             //                 Processador_data_master.address
		.Processador_data_master_waitrequest           (processador_data_master_waitrequest),                         //                                        .waitrequest
		.Processador_data_master_byteenable            (processador_data_master_byteenable),                          //                                        .byteenable
		.Processador_data_master_read                  (processador_data_master_read),                                //                                        .read
		.Processador_data_master_readdata              (processador_data_master_readdata),                            //                                        .readdata
		.Processador_data_master_write                 (processador_data_master_write),                               //                                        .write
		.Processador_data_master_writedata             (processador_data_master_writedata),                           //                                        .writedata
		.Processador_data_master_debugaccess           (processador_data_master_debugaccess),                         //                                        .debugaccess
		.Processador_instruction_master_address        (processador_instruction_master_address),                      //          Processador_instruction_master.address
		.Processador_instruction_master_waitrequest    (processador_instruction_master_waitrequest),                  //                                        .waitrequest
		.Processador_instruction_master_read           (processador_instruction_master_read),                         //                                        .read
		.Processador_instruction_master_readdata       (processador_instruction_master_readdata),                     //                                        .readdata
		.Conduit_Img_1_Escrita_write                   (mm_interconnect_0_conduit_img_1_escrita_write),               //                   Conduit_Img_1_Escrita.write
		.Conduit_Img_1_Escrita_writedata               (mm_interconnect_0_conduit_img_1_escrita_writedata),           //                                        .writedata
		.Conduit_Img_1_Leitura_read                    (mm_interconnect_0_conduit_img_1_leitura_read),                //                   Conduit_Img_1_Leitura.read
		.Conduit_Img_1_Leitura_readdata                (mm_interconnect_0_conduit_img_1_leitura_readdata),            //                                        .readdata
		.Conduit_Img_2_Escrita_write                   (mm_interconnect_0_conduit_img_2_escrita_write),               //                   Conduit_Img_2_Escrita.write
		.Conduit_Img_2_Escrita_writedata               (mm_interconnect_0_conduit_img_2_escrita_writedata),           //                                        .writedata
		.Conduit_Img_2_Leitura_read                    (mm_interconnect_0_conduit_img_2_leitura_read),                //                   Conduit_Img_2_Leitura.read
		.Conduit_Img_2_Leitura_readdata                (mm_interconnect_0_conduit_img_2_leitura_readdata),            //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.Medidor_Escrita_write                         (mm_interconnect_0_medidor_escrita_write),                     //                         Medidor_Escrita.write
		.Medidor_Escrita_writedata                     (mm_interconnect_0_medidor_escrita_writedata),                 //                                        .writedata
		.Medidor_Leitura_read                          (mm_interconnect_0_medidor_leitura_read),                      //                         Medidor_Leitura.read
		.Medidor_Leitura_readdata                      (mm_interconnect_0_medidor_leitura_readdata),                  //                                        .readdata
		.MemoriaImg1_s1_address                        (mm_interconnect_0_memoriaimg1_s1_address),                    //                          MemoriaImg1_s1.address
		.MemoriaImg1_s1_write                          (mm_interconnect_0_memoriaimg1_s1_write),                      //                                        .write
		.MemoriaImg1_s1_readdata                       (mm_interconnect_0_memoriaimg1_s1_readdata),                   //                                        .readdata
		.MemoriaImg1_s1_writedata                      (mm_interconnect_0_memoriaimg1_s1_writedata),                  //                                        .writedata
		.MemoriaImg1_s1_chipselect                     (mm_interconnect_0_memoriaimg1_s1_chipselect),                 //                                        .chipselect
		.MemoriaImg1_s1_clken                          (mm_interconnect_0_memoriaimg1_s1_clken),                      //                                        .clken
		.MemoriaImg1_s1_debugaccess                    (mm_interconnect_0_memoriaimg1_s1_debugaccess),                //                                        .debugaccess
		.MemoriaImg2_s1_address                        (mm_interconnect_0_memoriaimg2_s1_address),                    //                          MemoriaImg2_s1.address
		.MemoriaImg2_s1_write                          (mm_interconnect_0_memoriaimg2_s1_write),                      //                                        .write
		.MemoriaImg2_s1_readdata                       (mm_interconnect_0_memoriaimg2_s1_readdata),                   //                                        .readdata
		.MemoriaImg2_s1_writedata                      (mm_interconnect_0_memoriaimg2_s1_writedata),                  //                                        .writedata
		.MemoriaImg2_s1_chipselect                     (mm_interconnect_0_memoriaimg2_s1_chipselect),                 //                                        .chipselect
		.MemoriaImg2_s1_clken                          (mm_interconnect_0_memoriaimg2_s1_clken),                      //                                        .clken
		.MemoriaImg2_s1_debugaccess                    (mm_interconnect_0_memoriaimg2_s1_debugaccess),                //                                        .debugaccess
		.MemoriaPrograma_s1_address                    (mm_interconnect_0_memoriaprograma_s1_address),                //                      MemoriaPrograma_s1.address
		.MemoriaPrograma_s1_write                      (mm_interconnect_0_memoriaprograma_s1_write),                  //                                        .write
		.MemoriaPrograma_s1_readdata                   (mm_interconnect_0_memoriaprograma_s1_readdata),               //                                        .readdata
		.MemoriaPrograma_s1_writedata                  (mm_interconnect_0_memoriaprograma_s1_writedata),              //                                        .writedata
		.MemoriaPrograma_s1_byteenable                 (mm_interconnect_0_memoriaprograma_s1_byteenable),             //                                        .byteenable
		.MemoriaPrograma_s1_chipselect                 (mm_interconnect_0_memoriaprograma_s1_chipselect),             //                                        .chipselect
		.MemoriaPrograma_s1_clken                      (mm_interconnect_0_memoriaprograma_s1_clken),                  //                                        .clken
		.Processador_debug_mem_slave_address           (mm_interconnect_0_processador_debug_mem_slave_address),       //             Processador_debug_mem_slave.address
		.Processador_debug_mem_slave_write             (mm_interconnect_0_processador_debug_mem_slave_write),         //                                        .write
		.Processador_debug_mem_slave_read              (mm_interconnect_0_processador_debug_mem_slave_read),          //                                        .read
		.Processador_debug_mem_slave_readdata          (mm_interconnect_0_processador_debug_mem_slave_readdata),      //                                        .readdata
		.Processador_debug_mem_slave_writedata         (mm_interconnect_0_processador_debug_mem_slave_writedata),     //                                        .writedata
		.Processador_debug_mem_slave_byteenable        (mm_interconnect_0_processador_debug_mem_slave_byteenable),    //                                        .byteenable
		.Processador_debug_mem_slave_waitrequest       (mm_interconnect_0_processador_debug_mem_slave_waitrequest),   //                                        .waitrequest
		.Processador_debug_mem_slave_debugaccess       (mm_interconnect_0_processador_debug_mem_slave_debugaccess),   //                                        .debugaccess
		.Subtrator_Leitura_read                        (mm_interconnect_0_subtrator_leitura_read),                    //                       Subtrator_Leitura.read
		.Subtrator_Leitura_readdata                    (mm_interconnect_0_subtrator_leitura_readdata)                 //                                        .readdata
	);

	SistemaEmbarcado_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (processador_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                        // reset_in0.reset
		.reset_in1      (processador_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),        // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),    //          .reset_req
		.reset_req_in0  (1'b0),                                  // (terminated)
		.reset_req_in1  (1'b0),                                  // (terminated)
		.reset_in2      (1'b0),                                  // (terminated)
		.reset_req_in2  (1'b0),                                  // (terminated)
		.reset_in3      (1'b0),                                  // (terminated)
		.reset_req_in3  (1'b0),                                  // (terminated)
		.reset_in4      (1'b0),                                  // (terminated)
		.reset_req_in4  (1'b0),                                  // (terminated)
		.reset_in5      (1'b0),                                  // (terminated)
		.reset_req_in5  (1'b0),                                  // (terminated)
		.reset_in6      (1'b0),                                  // (terminated)
		.reset_req_in6  (1'b0),                                  // (terminated)
		.reset_in7      (1'b0),                                  // (terminated)
		.reset_req_in7  (1'b0),                                  // (terminated)
		.reset_in8      (1'b0),                                  // (terminated)
		.reset_req_in8  (1'b0),                                  // (terminated)
		.reset_in9      (1'b0),                                  // (terminated)
		.reset_req_in9  (1'b0),                                  // (terminated)
		.reset_in10     (1'b0),                                  // (terminated)
		.reset_req_in10 (1'b0),                                  // (terminated)
		.reset_in11     (1'b0),                                  // (terminated)
		.reset_req_in11 (1'b0),                                  // (terminated)
		.reset_in12     (1'b0),                                  // (terminated)
		.reset_req_in12 (1'b0),                                  // (terminated)
		.reset_in13     (1'b0),                                  // (terminated)
		.reset_req_in13 (1'b0),                                  // (terminated)
		.reset_in14     (1'b0),                                  // (terminated)
		.reset_req_in14 (1'b0),                                  // (terminated)
		.reset_in15     (1'b0),                                  // (terminated)
		.reset_req_in15 (1'b0)                                   // (terminated)
	);

endmodule
